`include "prefix.v"

module floatAdd(a, b, res, clk);
	dff(a, b, 3);
